module enemy_bit_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin

		if(({row_reg, col_reg}>=12'b000000000000) && ({row_reg, col_reg}<12'b000101011011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b000101011011)) color_data = 12'b110111101101;

		if(({row_reg, col_reg}>=12'b000101011100) && ({row_reg, col_reg}<12'b000110001101)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b000110001101)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b000110001110)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==12'b000110001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b000110010000)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b000110010001) && ({row_reg, col_reg}<12'b000110011001)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b000110011001)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b000110011010)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b000110011011)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b000110011100)) color_data = 12'b110111101101;

		if(({row_reg, col_reg}>=12'b000110011101) && ({row_reg, col_reg}<12'b000111001110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b000111001110)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b000111001111)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b000111010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b000111010001) && ({row_reg, col_reg}<12'b000111011001)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b000111011001)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b000111011010)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b000111011011)) color_data = 12'b101111001011;

		if(({row_reg, col_reg}>=12'b000111011100) && ({row_reg, col_reg}<12'b001000000111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001000000111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b001000001000) && ({row_reg, col_reg}<12'b001000001110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001000001110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001000001111)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b001000010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001000010001)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001000010010)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001000010011)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001000010100)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b001000010101)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001000010110)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b001000010111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001000011000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001000011001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b001000011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001000011011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b001000011100) && ({row_reg, col_reg}<12'b001000100011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001000100011)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b001000100100) && ({row_reg, col_reg}<12'b001001000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001001000110)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b001001000111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}>=12'b001001001000) && ({row_reg, col_reg}<12'b001001001111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001001001111)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b001001010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001001010001)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001001010010)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001001010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001001010101)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==12'b001001010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001001010111)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==12'b001001011000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001001011001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b001001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001001011011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b001001011100) && ({row_reg, col_reg}<12'b001001100010)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001001100010)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b001001100011)) color_data = 12'b101111001011;

		if(({row_reg, col_reg}>=12'b001001100100) && ({row_reg, col_reg}<12'b001010000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001010000110)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b001010000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001010001000)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=12'b001010001001) && ({row_reg, col_reg}<12'b001010001110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001010001110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001010001111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b001010010000)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==12'b001010010001)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001010010010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b001010010011)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b001010010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001010010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b001010010110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b001010010111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001010011000)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001010011001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b001010011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001010011011)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b001010011100) && ({row_reg, col_reg}<12'b001010100001)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001010100001)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b001010100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001010100011)) color_data = 12'b101110111010;

		if(({row_reg, col_reg}>=12'b001010100100) && ({row_reg, col_reg}<12'b001011000111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001011000111)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b001011001000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001011001001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=12'b001011001010) && ({row_reg, col_reg}<12'b001011001100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}>=12'b001011001100) && ({row_reg, col_reg}<12'b001011001110)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001011001110)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==12'b001011001111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001011010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001011010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001011010010)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b001011010011)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==12'b001011010100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b001011010101)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b001011010110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b001011010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b001011011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001011011001)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b001011011010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001011011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001011011100)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}>=12'b001011011101) && ({row_reg, col_reg}<12'b001011011111)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001011011111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001011100000)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b001011100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001011100010)) color_data = 12'b101110111010;

		if(({row_reg, col_reg}>=12'b001011100011) && ({row_reg, col_reg}<12'b001100001000)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001100001000)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b001100001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001100001010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b001100001011)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==12'b001100001100)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b001100001101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001100001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001100001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001100010000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001100010001)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b001100010010)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==12'b001100010011)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}>=12'b001100010100) && ({row_reg, col_reg}<12'b001100010110)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==12'b001100010110)) color_data = 12'b011000110100;
		if(({row_reg, col_reg}==12'b001100010111)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b001100011000)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==12'b001100011001)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b001100011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b001100011011) && ({row_reg, col_reg}<12'b001100011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001100011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b001100011110)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b001100011111)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b001100100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b001100100001)) color_data = 12'b101010111010;

		if(({row_reg, col_reg}>=12'b001100100010) && ({row_reg, col_reg}<12'b001101001000)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001101001000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001101001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001101001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001101001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001101001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001101001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001101001110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b001101001111)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b001101010000)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b001101010001)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b001101010010)) color_data = 12'b011001000101;
		if(({row_reg, col_reg}==12'b001101010011)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}>=12'b001101010100) && ({row_reg, col_reg}<12'b001101010111)) color_data = 12'b101101100100;
		if(({row_reg, col_reg}==12'b001101010111)) color_data = 12'b100101010100;
		if(({row_reg, col_reg}==12'b001101011000)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}==12'b001101011001)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b001101011010)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b001101011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001101011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001101011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001101011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001101011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001101100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001101100001)) color_data = 12'b110111011100;

		if(({row_reg, col_reg}>=12'b001101100010) && ({row_reg, col_reg}<12'b001110001000)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001110001000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001110001001)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}>=12'b001110001010) && ({row_reg, col_reg}<12'b001110001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001110001100)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b001110001101)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==12'b001110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001110001111)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==12'b001110010000)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}==12'b001110010001)) color_data = 12'b010001001000;
		if(({row_reg, col_reg}==12'b001110010010)) color_data = 12'b010101011000;
		if(({row_reg, col_reg}==12'b001110010011)) color_data = 12'b101001100111;
		if(({row_reg, col_reg}==12'b001110010100)) color_data = 12'b110010000101;
		if(({row_reg, col_reg}==12'b001110010101)) color_data = 12'b110010010110;
		if(({row_reg, col_reg}==12'b001110010110)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}==12'b001110010111)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}==12'b001110011000)) color_data = 12'b010001011000;
		if(({row_reg, col_reg}==12'b001110011001)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}==12'b001110011010)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b001110011011)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b001110011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001110011101)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b001110011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001110011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001110100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001110100001)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b001110100010) && ({row_reg, col_reg}<12'b001111000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001111000110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b001111000111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b001111001000)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==12'b001111001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001111001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b001111001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001111001100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b001111001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001111001110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b001111001111)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b001111010000)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}==12'b001111010001)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b001111010010)) color_data = 12'b010101101011;
		if(({row_reg, col_reg}==12'b001111010011)) color_data = 12'b011001111011;
		if(({row_reg, col_reg}==12'b001111010100)) color_data = 12'b101001110111;
		if(({row_reg, col_reg}==12'b001111010101)) color_data = 12'b110001110100;
		if(({row_reg, col_reg}==12'b001111010110)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==12'b001111010111)) color_data = 12'b011001111100;
		if(({row_reg, col_reg}==12'b001111011000)) color_data = 12'b010001011010;
		if(({row_reg, col_reg}==12'b001111011001)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b001111011010)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}==12'b001111011011)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==12'b001111011100)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b001111011101)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}>=12'b001111011110) && ({row_reg, col_reg}<12'b001111100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b001111100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b001111100001)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b001111100010)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b001111100011) && ({row_reg, col_reg}<12'b001111100101)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b001111100101) && ({row_reg, col_reg}<12'b010000000100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010000000100)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b010000000101)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b010000000110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b010000000111)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==12'b010000001000)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b010000001001)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010000001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010000001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010000001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010000001101)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b010000001110)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b010000001111)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010000010000)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}>=12'b010000010001) && ({row_reg, col_reg}<12'b010000010011)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b010000010011)) color_data = 12'b011101101010;
		if(({row_reg, col_reg}==12'b010000010100)) color_data = 12'b101101110101;
		if(({row_reg, col_reg}==12'b010000010101)) color_data = 12'b110001110100;
		if(({row_reg, col_reg}==12'b010000010110)) color_data = 12'b100101101000;
		if(({row_reg, col_reg}==12'b010000010111)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==12'b010000011000)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}==12'b010000011001)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}>=12'b010000011010) && ({row_reg, col_reg}<12'b010000011100)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010000011100)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b010000011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010000011110)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b010000011111)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b010000100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010000100001)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b010000100010)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b010000100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b010000100100)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b010000100101)) color_data = 12'b110111101101;

		if(({row_reg, col_reg}>=12'b010000100110) && ({row_reg, col_reg}<12'b010001000011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010001000011)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b010001000100)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b010001000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010001000110)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b010001000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010001001000)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b010001001001)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b010001001010)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b010001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010001001100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==12'b010001001101)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}>=12'b010001001110) && ({row_reg, col_reg}<12'b010001010001)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010001010001)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}==12'b010001010010)) color_data = 12'b010101011000;
		if(({row_reg, col_reg}==12'b010001010011)) color_data = 12'b101001010101;
		if(({row_reg, col_reg}==12'b010001010100)) color_data = 12'b110001100100;
		if(({row_reg, col_reg}==12'b010001010101)) color_data = 12'b101101100100;
		if(({row_reg, col_reg}==12'b010001010110)) color_data = 12'b101101010100;
		if(({row_reg, col_reg}==12'b010001010111)) color_data = 12'b100001000110;
		if(({row_reg, col_reg}==12'b010001011000)) color_data = 12'b010001011000;
		if(({row_reg, col_reg}==12'b010001011001)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}>=12'b010001011010) && ({row_reg, col_reg}<12'b010001011100)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010001011100)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b010001011101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==12'b010001011110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010001011111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b010001100000)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010001100001)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b010001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010001100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010001100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010001100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010001100110)) color_data = 12'b110011001011;

		if(({row_reg, col_reg}==12'b010001100111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b010010000000) && ({row_reg, col_reg}<12'b010010000011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010010000011)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b010010000100)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b010010000101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010010000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010010000111)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}>=12'b010010001000) && ({row_reg, col_reg}<12'b010010001011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b010010001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010010001100)) color_data = 12'b000000000001;
		if(({row_reg, col_reg}==12'b010010001101)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}>=12'b010010001110) && ({row_reg, col_reg}<12'b010010010010)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010010010010)) color_data = 12'b100001000101;
		if(({row_reg, col_reg}==12'b010010010011)) color_data = 12'b011101000101;
		if(({row_reg, col_reg}==12'b010010010100)) color_data = 12'b011001011000;
		if(({row_reg, col_reg}==12'b010010010101)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}==12'b010010010110)) color_data = 12'b011101010111;
		if(({row_reg, col_reg}==12'b010010010111)) color_data = 12'b100001000100;
		if(({row_reg, col_reg}==12'b010010011000)) color_data = 12'b011001000110;
		if(({row_reg, col_reg}>=12'b010010011001) && ({row_reg, col_reg}<12'b010010011100)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010010011100)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b010010011101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==12'b010010011110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010010011111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}>=12'b010010100000) && ({row_reg, col_reg}<12'b010010100010)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b010010100010)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010010100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010010100101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==12'b010010100110)) color_data = 12'b100110101001;

		if(({row_reg, col_reg}==12'b010010100111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b010011000000) && ({row_reg, col_reg}<12'b010011000011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010011000011)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b010011000100)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b010011000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010011000110)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010011000111)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010011001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010011001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010011001010)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b010011001011)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b010011001100)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010011001101)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010011001110)) color_data = 12'b001100110101;
		if(({row_reg, col_reg}>=12'b010011001111) && ({row_reg, col_reg}<12'b010011010010)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010011010010)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}>=12'b010011010011) && ({row_reg, col_reg}<12'b010011010101)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010011010101)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}>=12'b010011010110) && ({row_reg, col_reg}<12'b010011011000)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010011011000)) color_data = 12'b010000110101;
		if(({row_reg, col_reg}>=12'b010011011001) && ({row_reg, col_reg}<12'b010011011100)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010011011100)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b010011011101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==12'b010011011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010011011111)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b010011100000)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b010011100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010011100011)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b010011100100)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010011100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010011100110)) color_data = 12'b110011001011;

		if(({row_reg, col_reg}==12'b010011100111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b010100000000) && ({row_reg, col_reg}<12'b010100000100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010100000100)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b010100000101)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b010100000110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b010100000111)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b010100001000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010100001001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010100001010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010100001011)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b010100001100)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b010100001101)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010100001110)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}>=12'b010100001111) && ({row_reg, col_reg}<12'b010100010010)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010100010010)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}>=12'b010100010011) && ({row_reg, col_reg}<12'b010100011000)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b010100011000)) color_data = 12'b001100110101;
		if(({row_reg, col_reg}>=12'b010100011001) && ({row_reg, col_reg}<12'b010100011011)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010100011011)) color_data = 12'b001100110101;
		if(({row_reg, col_reg}==12'b010100011100)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b010100011101)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==12'b010100011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010100011111)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b010100100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010100100001)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010100100010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b010100100011)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==12'b010100100100)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b010100100101)) color_data = 12'b110111101101;

		if(({row_reg, col_reg}>=12'b010100100110) && ({row_reg, col_reg}<12'b010101000111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010101000111)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b010101001000)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b010101001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010101001010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010101001011)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010101001100)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==12'b010101001101)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==12'b010101001110)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}>=12'b010101001111) && ({row_reg, col_reg}<12'b010101010001)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b010101010001)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==12'b010101010010)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010101010011)) color_data = 12'b001000010011;
		if(({row_reg, col_reg}==12'b010101010100)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==12'b010101010101)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b010101010110)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}>=12'b010101010111) && ({row_reg, col_reg}<12'b010101011001)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010101011001)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b010101011010)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b010101011011)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b010101011100)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==12'b010101011101)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==12'b010101011110)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==12'b010101011111)) color_data = 12'b001000100010;
		if(({row_reg, col_reg}==12'b010101100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010101100001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=12'b010101100010) && ({row_reg, col_reg}<12'b010101100100)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b010101100100)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b010101100101) && ({row_reg, col_reg}<12'b010110001000)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}>=12'b010110001000) && ({row_reg, col_reg}<12'b010110001010)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b010110001010)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==12'b010110001011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b010110001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010110001101)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b010110001110)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010110001111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==12'b010110010000)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010110010001)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b010110010010)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b010110010011)) color_data = 12'b001101000111;
		if(({row_reg, col_reg}>=12'b010110010100) && ({row_reg, col_reg}<12'b010110010110)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b010110010110)) color_data = 12'b010001011000;
		if(({row_reg, col_reg}==12'b010110010111)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010110011000)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==12'b010110011001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}>=12'b010110011010) && ({row_reg, col_reg}<12'b010110011100)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010110011100)) color_data = 12'b000100010010;
		if(({row_reg, col_reg}==12'b010110011101)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==12'b010110011110)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b010110011111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b010110100000)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b010110100001)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b010110100010) && ({row_reg, col_reg}<12'b010111000111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b010111000111)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b010111001000)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}>=12'b010111001001) && ({row_reg, col_reg}<12'b010111001011)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b010111001011)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b010111001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010111001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b010111001110)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==12'b010111001111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b010111010000)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b010111010001)) color_data = 12'b001100110101;
		if(({row_reg, col_reg}==12'b010111010010)) color_data = 12'b001101000111;
		if(({row_reg, col_reg}==12'b010111010011)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b010111010100)) color_data = 12'b010001011010;
		if(({row_reg, col_reg}==12'b010111010101)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}>=12'b010111010110) && ({row_reg, col_reg}<12'b010111011000)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b010111011000)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b010111011001)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==12'b010111011010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==12'b010111011011)) color_data = 12'b000100000001;
		if(({row_reg, col_reg}==12'b010111011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==12'b010111011101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b010111011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111011111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b010111100000)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b010111100001)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b010111100010)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b010111100011) && ({row_reg, col_reg}<12'b011000000111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011000000111)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011000001000)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b011000001001)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b011000001010)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011000001011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000001100)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b011000001101)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b011000001110)) color_data = 12'b001000010001;
		if(({row_reg, col_reg}==12'b011000001111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==12'b011000010000)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b011000010001)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b011000010010)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}==12'b011000010011)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}>=12'b011000010100) && ({row_reg, col_reg}<12'b011000010110)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}>=12'b011000010110) && ({row_reg, col_reg}<12'b011000011000)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b011000011000)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}==12'b011000011001)) color_data = 12'b001100100101;
		if(({row_reg, col_reg}==12'b011000011010)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==12'b011000011011)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==12'b011000011100)) color_data = 12'b000100010001;
		if(({row_reg, col_reg}==12'b011000011101)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}>=12'b011000011110) && ({row_reg, col_reg}<12'b011000100000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000100000)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b011000100001)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011000100010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011000100011)) color_data = 12'b110111101101;

		if(({row_reg, col_reg}>=12'b011000100100) && ({row_reg, col_reg}<12'b011001000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011001000110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011001000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011001001000)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b011001001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011001001010)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011001001011)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011001001100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b011001001101)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b011001001110)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==12'b011001001111)) color_data = 12'b101101110100;
		if(({row_reg, col_reg}==12'b011001010000)) color_data = 12'b011001000011;
		if(({row_reg, col_reg}==12'b011001010001)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b011001010010)) color_data = 12'b001000100110;
		if(({row_reg, col_reg}==12'b011001010011)) color_data = 12'b001101001000;
		if(({row_reg, col_reg}>=12'b011001010100) && ({row_reg, col_reg}<12'b011001010111)) color_data = 12'b010001011001;
		if(({row_reg, col_reg}==12'b011001010111)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}==12'b011001011000)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b011001011001)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b011001011010)) color_data = 12'b100101100100;
		if(({row_reg, col_reg}==12'b011001011011)) color_data = 12'b101001010100;
		if(({row_reg, col_reg}==12'b011001011100)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==12'b011001011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011001011110)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b011001011111)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==12'b011001100000)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b011001100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011001100010)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b011001100011)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011001100100)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b011001100101) && ({row_reg, col_reg}<12'b011010000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011010000110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011010000111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b011010001000)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b011010001001)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011010001010)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b011010001011)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011010001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011010001101)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}>=12'b011010001110) && ({row_reg, col_reg}<12'b011010010000)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==12'b011010010000)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==12'b011010010001)) color_data = 12'b001100100010;
		if(({row_reg, col_reg}==12'b011010010010)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==12'b011010010011)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b011010010100)) color_data = 12'b001100110111;
		if(({row_reg, col_reg}==12'b011010010101)) color_data = 12'b001101000111;
		if(({row_reg, col_reg}==12'b011010010110)) color_data = 12'b001100110110;
		if(({row_reg, col_reg}==12'b011010010111)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==12'b011010011000)) color_data = 12'b010000100011;
		if(({row_reg, col_reg}==12'b011010011001)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==12'b011010011010)) color_data = 12'b011101000011;
		if(({row_reg, col_reg}==12'b011010011011)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==12'b011010011100)) color_data = 12'b011101000100;
		if(({row_reg, col_reg}==12'b011010011101)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011010011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011010011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011010100000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011010100001)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011010100010)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b011010100011)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011010100100)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b011010100101) && ({row_reg, col_reg}<12'b011011000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011011000110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011011000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011001000)) color_data = 12'b010000110100;
		if(({row_reg, col_reg}==12'b011011001001)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b011011001010)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b011011001011)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b011011001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b011011001101)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011011001110)) color_data = 12'b010101000100;
		if(({row_reg, col_reg}==12'b011011001111)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==12'b011011010000)) color_data = 12'b010000010010;
		if(({row_reg, col_reg}==12'b011011010001)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==12'b011011010010)) color_data = 12'b110010000100;
		if(({row_reg, col_reg}==12'b011011010011)) color_data = 12'b100001100011;
		if(({row_reg, col_reg}==12'b011011010100)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==12'b011011010101)) color_data = 12'b001000100110;
		if(({row_reg, col_reg}==12'b011011010110)) color_data = 12'b010000110011;
		if(({row_reg, col_reg}==12'b011011010111)) color_data = 12'b101110000100;
		if(({row_reg, col_reg}==12'b011011011000)) color_data = 12'b110001100100;
		if(({row_reg, col_reg}==12'b011011011001)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==12'b011011011010)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==12'b011011011011)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==12'b011011011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011011101)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011011011110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011011011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011011100000)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011011100001)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011011100010)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b011011100011)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011011100100)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b011011100101) && ({row_reg, col_reg}<12'b011100000111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011100000111)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011100001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011100001001)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b011100001010)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011100001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011100001100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011100001101)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b011100001110)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011100001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b011100010000)) color_data = 12'b010000100010;
		if(({row_reg, col_reg}==12'b011100010001)) color_data = 12'b110001010100;
		if(({row_reg, col_reg}==12'b011100010010)) color_data = 12'b101101010100;
		if(({row_reg, col_reg}==12'b011100010011)) color_data = 12'b100101010011;
		if(({row_reg, col_reg}==12'b011100010100)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b011100010101)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==12'b011100010110)) color_data = 12'b010100110011;
		if(({row_reg, col_reg}==12'b011100010111)) color_data = 12'b101001100100;
		if(({row_reg, col_reg}==12'b011100011000)) color_data = 12'b110001010100;
		if(({row_reg, col_reg}==12'b011100011001)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==12'b011100011010)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b011100011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011100011100)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011100011101)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b011100011110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011100011111)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b011100100000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011100100001)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011100100010)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b011100100011) && ({row_reg, col_reg}<12'b011101000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011101000110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011101000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b011101001000)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011101001001)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b011101001010)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011101001011)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011101001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011101001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011101001110)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b011101001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011101010000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011101010001)) color_data = 12'b100101000100;
		if(({row_reg, col_reg}==12'b011101010010)) color_data = 12'b100100110100;
		if(({row_reg, col_reg}==12'b011101010011)) color_data = 12'b010100100011;
		if(({row_reg, col_reg}>=12'b011101010100) && ({row_reg, col_reg}<12'b011101010111)) color_data = 12'b001100010010;
		if(({row_reg, col_reg}==12'b011101010111)) color_data = 12'b011100110011;
		if(({row_reg, col_reg}==12'b011101011000)) color_data = 12'b101001000100;
		if(({row_reg, col_reg}==12'b011101011001)) color_data = 12'b100001010101;
		if(({row_reg, col_reg}==12'b011101011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011101011011)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011101011100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011101011101)) color_data = 12'b010101000101;
		if(({row_reg, col_reg}==12'b011101011110)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}>=12'b011101011111) && ({row_reg, col_reg}<12'b011101100001)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011101100001)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011101100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011101100011)) color_data = 12'b110111011100;

		if(({row_reg, col_reg}>=12'b011101100100) && ({row_reg, col_reg}<12'b011110000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011110000110)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}==12'b011110000111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011110001000)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b011110001001)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}>=12'b011110001010) && ({row_reg, col_reg}<12'b011110001100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011110001100)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011110001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011110001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011110001111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011110010000)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011110010001)) color_data = 12'b011001010110;
		if(({row_reg, col_reg}==12'b011110010010)) color_data = 12'b001100010011;
		if(({row_reg, col_reg}==12'b011110010011)) color_data = 12'b001100100100;
		if(({row_reg, col_reg}==12'b011110010100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011110010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011110010110)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b011110010111)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b011110011000)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b011110011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b011110011010)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011110011011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011110011100)) color_data = 12'b001100100011;
		if(({row_reg, col_reg}==12'b011110011101)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==12'b011110011110)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011110011111)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011110100000)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011110100001)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011110100010)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b011110100011)) color_data = 12'b101010101001;

		if(({row_reg, col_reg}>=12'b011110100100) && ({row_reg, col_reg}<12'b011111000110)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011111000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011111000111)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b011111001000)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b011111001001)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b011111001010) && ({row_reg, col_reg}<12'b011111001100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011111001100)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b011111001101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b011111001110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b011111001111)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011111010000)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011111010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011111010010)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b011111010011)) color_data = 12'b001100110101;
		if(({row_reg, col_reg}==12'b011111010100)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b011111010101)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b011111010110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==12'b011111010111)) color_data = 12'b001000100101;
		if(({row_reg, col_reg}==12'b011111011000)) color_data = 12'b001100110101;
		if(({row_reg, col_reg}==12'b011111011001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b011111011010)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}>=12'b011111011011) && ({row_reg, col_reg}<12'b011111011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011111011101)) color_data = 12'b110111101100;
		if(({row_reg, col_reg}>=12'b011111011110) && ({row_reg, col_reg}<12'b011111100001)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b011111100001)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b011111100010)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b011111100011)) color_data = 12'b001000100011;
		if(({row_reg, col_reg}==12'b011111100100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b011111100101)) color_data = 12'b111011111101;

		if(({row_reg, col_reg}>=12'b011111100110) && ({row_reg, col_reg}<12'b100000000101)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100000000101)) color_data = 12'b101111001011;
		if(({row_reg, col_reg}==12'b100000000110)) color_data = 12'b010001000100;
		if(({row_reg, col_reg}==12'b100000000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100000001000)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b100000001001) && ({row_reg, col_reg}<12'b100000001101)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100000001101)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100000001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100000001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b100000010000)) color_data = 12'b110011011011;
		if(({row_reg, col_reg}==12'b100000010001)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100000010010)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b100000010011)) color_data = 12'b001000100100;
		if(({row_reg, col_reg}==12'b100000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100000010101)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}>=12'b100000010110) && ({row_reg, col_reg}<12'b100000011000)) color_data = 12'b001100110101;
		if(({row_reg, col_reg}==12'b100000011000)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==12'b100000011001)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b100000011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100000011011)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b100000011100)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100000011101)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b100000011110) && ({row_reg, col_reg}<12'b100000100001)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100000100001)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100000100010)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100000100011)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100000100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100000100101)) color_data = 12'b110111101101;

		if(({row_reg, col_reg}>=12'b100000100110) && ({row_reg, col_reg}<12'b100001000011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100001000011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100001000100)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100001000101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001000110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100001000111)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b100001001000) && ({row_reg, col_reg}<12'b100001001101)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100001001101)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b100001001110)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001001111)) color_data = 12'b001100110011;
		if(({row_reg, col_reg}==12'b100001010000)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100001010001)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100001010010)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100001010011)) color_data = 12'b010101010110;
		if(({row_reg, col_reg}==12'b100001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100001010101)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==12'b100001010110)) color_data = 12'b010001000101;
		if(({row_reg, col_reg}==12'b100001010111)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==12'b100001011000)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b100001011001)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100001011011)) color_data = 12'b001000010010;
		if(({row_reg, col_reg}==12'b100001011100)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b100001011101)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}>=12'b100001011110) && ({row_reg, col_reg}<12'b100001100010)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100001100010)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100001100011)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100001100100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100001100101)) color_data = 12'b100010001000;

		if(({row_reg, col_reg}>=12'b100001100110) && ({row_reg, col_reg}<12'b100010000100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100010000100)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100010000101)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b100010000110)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b100010000111) && ({row_reg, col_reg}<12'b100010001101)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b100010001110)) color_data = 12'b001100110100;
		if(({row_reg, col_reg}==12'b100010001111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=12'b100010010000) && ({row_reg, col_reg}<12'b100010010011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}>=12'b100010010011) && ({row_reg, col_reg}<12'b100010010101)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b100010010101)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b100010010110)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}==12'b100010010111)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}>=12'b100010011000) && ({row_reg, col_reg}<12'b100010011010)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100010011010)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b100010011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100010011100)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100010011101)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}>=12'b100010011110) && ({row_reg, col_reg}<12'b100010100011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100010100011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100010100100)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==12'b100010100101)) color_data = 12'b100110101001;

		if(({row_reg, col_reg}>=12'b100010100110) && ({row_reg, col_reg}<12'b100011001011)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100011001011)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100011001100)) color_data = 12'b110011001011;
		if(({row_reg, col_reg}==12'b100011001101)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}==12'b100011001110)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}>=12'b100011001111) && ({row_reg, col_reg}<12'b100011011010)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100011011010)) color_data = 12'b111011111101;
		if(({row_reg, col_reg}==12'b100011011011)) color_data = 12'b110111011100;
		if(({row_reg, col_reg}==12'b100011011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100011011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b100011011110)) color_data = 12'b110111101101;

		if(({row_reg, col_reg}>=12'b100011011111) && ({row_reg, col_reg}<12'b100100001100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100100001100)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b100100001101)) color_data = 12'b110011011100;
		if(({row_reg, col_reg}>=12'b100100001110) && ({row_reg, col_reg}<12'b100100011100)) color_data = 12'b111011101101;
		if(({row_reg, col_reg}==12'b100100011100)) color_data = 12'b110111101101;
		if(({row_reg, col_reg}==12'b100100011101)) color_data = 12'b110111011100;




		if(({row_reg, col_reg}>=12'b100100011110) && ({row_reg, col_reg}<=12'b100111100111)) color_data = 12'b111011101101;
	end
endmodule